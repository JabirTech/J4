module Adder(A, B);

input [3:0] A, B;
output C;

assign C = A + B; 

endmodule
