module NOTer(A); 

input [3:0] A; 
output C; 

assign C = ~A; 

endmodule
